--==============================================================================
--== Logisim goes FPGA automatic generated VHDL code                          ==
--==                                                                          ==
--==                                                                          ==
--== Project   : golden                                                       ==
--== Component : toplevel                                                     ==
--==                                                                          ==
--==============================================================================


LIBRARY ieee;
USE ieee.std_logic_1164.all;
USE ieee.numeric_std.all;

ENTITY toplevel IS
   PORT ( Clock_0                   : IN  std_logic;
          n_Block_die_1_0           : IN  std_logic;
          n_Block_die_2_0           : IN  std_logic;
          n_Block_die_3_0           : IN  std_logic;
          n_Block_die_4_0           : IN  std_logic;
          n_Mode_0                  : IN  std_logic;
          n_Reset_0                 : IN  std_logic;
          L1_0                      : OUT std_logic;
          L2_0                      : OUT std_logic;
          L3_0                      : OUT std_logic;
          L4_0                      : OUT std_logic;
          L5_0                      : OUT std_logic;
          L6_0                      : OUT std_logic;
          die1_DecimalPoint         : OUT std_logic;
          die1_Segment_A            : OUT std_logic;
          die1_Segment_B            : OUT std_logic;
          die1_Segment_C            : OUT std_logic;
          die1_Segment_D            : OUT std_logic;
          die1_Segment_E            : OUT std_logic;
          die1_Segment_F            : OUT std_logic;
          die1_Segment_G            : OUT std_logic;
          die2_DecimalPoint         : OUT std_logic;
          die2_Segment_A            : OUT std_logic;
          die2_Segment_B            : OUT std_logic;
          die2_Segment_C            : OUT std_logic;
          die2_Segment_D            : OUT std_logic;
          die2_Segment_E            : OUT std_logic;
          die2_Segment_F            : OUT std_logic;
          die2_Segment_G            : OUT std_logic;
          die3_DecimalPoint         : OUT std_logic;
          die3_Segment_A            : OUT std_logic;
          die3_Segment_B            : OUT std_logic;
          die3_Segment_C            : OUT std_logic;
          die3_Segment_D            : OUT std_logic;
          die3_Segment_E            : OUT std_logic;
          die3_Segment_F            : OUT std_logic;
          die3_Segment_G            : OUT std_logic;
          die4_DecimalPoint         : OUT std_logic;
          die4_Segment_A            : OUT std_logic;
          die4_Segment_B            : OUT std_logic;
          die4_Segment_C            : OUT std_logic;
          die4_Segment_D            : OUT std_logic;
          die4_Segment_E            : OUT std_logic;
          die4_Segment_F            : OUT std_logic;
          die4_Segment_G            : OUT std_logic);
END toplevel;

